module asn1
