module main 

