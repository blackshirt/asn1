module main 


fn main() {
	// Basically this is a Kerberos PrincipalName data you sent to me
	const data = [u8(0x30), 0x15, 0xa0, 0x03, 0x02, 0x01, 0x01, 0xa1, 0x0e, 0x30, 0x0c, 0x1b, 0x0a,
	0x62, 0x6f, 0x62, 0x62, 0x61, 0x2d, 0x66, 0x65, 0x74, 0x74]
	p := PrincipalName{
		name_type: asn1.Int64.from_i64(1)
		name_string: [KerberosString.from_string('bobba-fett')!]
	}
	mut out := []u8{}
	p.encode(mut out)!
	assert out == data // should assert to true
}
